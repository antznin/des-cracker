ahmeda@makalu.15390:1556863729